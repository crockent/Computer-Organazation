--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:41:06 04/14/2024
-- Design Name:   
-- Module Name:   /home/manos/Documents/organosh/EX1V1/ALU_ex_test.vhd
-- Project Name:  EX1V1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: ALU_ex
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY ALU_ex_test IS
END ALU_ex_test;
 
ARCHITECTURE behavior OF ALU_ex_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT ALU_ex
    PORT(
         RF_A : IN  std_logic_vector(31 downto 0);
         RF_B : IN  std_logic_vector(31 downto 0);
         Immed : IN  std_logic_vector(31 downto 0);
         ALU_Bin_sel : IN  std_logic;
         ALU_Func : IN  std_logic_vector(3 downto 0);
         ALU_out : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal RF_A : std_logic_vector(31 downto 0) := (others => '0');
   signal RF_B : std_logic_vector(31 downto 0) := (others => '0');
   signal Immed : std_logic_vector(31 downto 0) := (others => '0');
   signal ALU_Bin_sel : std_logic := '0';
   signal ALU_Func : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal ALU_out : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
--   constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: ALU_ex PORT MAP (
          RF_A => RF_A,
          RF_B => RF_B,
          Immed => Immed,
          ALU_Bin_sel => ALU_Bin_sel,
          ALU_Func => ALU_Func,
          ALU_out => ALU_out
        );

--   -- Clock process definitions
--   <clock>_process :process
--   begin
--		<clock> <= '0';
--		wait for <clock>_period/2;
--		<clock> <= '1';
--		wait for <clock>_period/2;
--   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		RF_A <= x"00000001";
		RF_B <= x"00000002";
		ALU_Bin_sel<= '0';
		ALU_Func<="0000";
      wait for 100 ns;
		RF_A <= x"00000001";
		RF_B <= x"00000002";
		Immed <= x"00000003";
		ALU_Bin_sel<= '1';
		ALU_Func<="0000";
      wait for 100 ns;
		RF_A <= x"00000002";
		RF_B <= x"00000001";
		ALU_Bin_sel<= '0';
		ALU_Func<="0001";
      wait for 100 ns;
		RF_A <= x"00000002";
		RF_B <= x"00000001";
		ALU_Bin_sel<= '0';
		ALU_Func<="0010";
      wait for 100 ns;
		RF_A <= x"00000001";
		RF_B <= x"00000001";
		ALU_Bin_sel<= '0';
		ALU_Func<="0010";
      wait for 100 ns;
		RF_A <= x"00000002";
		RF_B <= x"00000001";
		ALU_Bin_sel<= '0';
		ALU_Func<="0011";
      wait for 100 ns;
		RF_A <= x"00000001";
		RF_B <= x"00000001";
		ALU_Bin_sel<= '0';
		ALU_Func<="0011";
      wait for 100 ns;
		RF_A <= x"00000002";
		RF_B <= x"00000001";
		ALU_Bin_sel<= '0';
		ALU_Func<="0100";
      wait for 100 ns;
		RF_A <= x"F0000002";
		RF_B <= x"00000001";
		ALU_Bin_sel<= '0';
		ALU_Func<="1000";
      wait for 100 ns;
		RF_A <= x"F000000F";
		ALU_Func<="1001";
      wait for 100 ns;
		RF_A <= x"F000000F";
		ALU_Func<="1010";
      wait for 100 ns;
		RF_A <= x"F000000F";
		ALU_Func<="1100";
      wait for 100 ns;
		RF_A <= x"F000000F";
		ALU_Func<="1101";
      wait for 100 ns;

      -- insert stimulus here 

      wait;
   end process;

END;
